
module INC_CTRL (
	probe);	

	input	[31:0]	probe;
endmodule
